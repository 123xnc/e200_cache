module mem(input           	   clk, we,
            input  [31:0]        a,
            input  [127:0]       wd,
            output [127:0]       rd);

  reg  [127:0] RAM[1023:0];

  assign rd = RAM[a[13:4]]; // set aligned

  integer i;
    
  initial begin
      for(i = 0; i <=1023; i=i+1) begin
        if(i == 0) RAM[i] = 128'h00C0006F063006132900081300000513;
                    //RAM[i] = 128'h00C0006F009006131280081300000513;
        else if (i == 1) RAM[i] = 128'h40B806B30025159302C50A6300150513;
        else if (i == 2) RAM[i] = 128'hFED702E30047071300C0006F10400713;
        else if (i == 3) RAM[i] = 128'hFEB72E23FEF5D8E300072583FFC72783;
        else if (i == 4) RAM[i] = 128'h0000806700000513FE5FF06F00F72023;

        else if (i == 16) RAM[i] = 128'h00000063000000790000000800000054;
        else if (i == 17) RAM[i] = 128'h00000037000000160000008300000081;
        else if (i == 18) RAM[i] = 128'h00000056000000140000002500000066;
        else if (i == 19) RAM[i] = 128'h00000090000000190000009800000074;
        else if (i == 20) RAM[i] = 128'h00000034000000180000007200000075;

        else if (i == 21) RAM[i] = 128'h00000043000000820000004900000005;
        else if (i == 22) RAM[i] = 128'h00000051000000210000004100000093;
        else if (i == 23) RAM[i] = 128'h00000039000000860000005800000088;
        else if (i == 24) RAM[i] = 128'h00000060000000270000008900000047;
        else if (i == 25) RAM[i] = 128'h00000067000000040000002000000094;

        else if (i == 26) RAM[i] = 128'h00000042000000690000008500000024;
        else if (i == 27) RAM[i] = 128'h00000077000000780000000300000022;
        else if (i == 28) RAM[i] = 128'h00000002000000760000007300000010;
        else if (i == 29) RAM[i] = 128'h00000100000000360000005500000045;
        else if (i == 30) RAM[i] = 128'h00000087000000170000004800000040;

        else if (i == 31) RAM[i] = 128'h00000015000000590000000700000062;
        else if (i == 32) RAM[i] = 128'h00000091000000280000006400000053;
        else if (i == 33) RAM[i] = 128'h00000095000000440000009200000009;
        else if (i == 34) RAM[i] = 128'h00000029000000680000003100000097;
        else if (i == 35) RAM[i] = 128'h00000035000000260000003300000012;

        else if (i == 36) RAM[i] = 128'h00000001000000130000005700000080;
        else if (i == 37) RAM[i] = 128'h00000023000000380000001100000052;
        else if (i == 38) RAM[i] = 128'h00000096000000060000005000000030;
        else if (i == 39) RAM[i] = 128'h00000061000000700000006500000099;
        else if (i == 40) RAM[i] = 128'h00000084000000710000004600000032;

	      else RAM[i] = 128'b0;
        // RAM[i] = 128'h00000013000000130000001300000013;
      end

      // RAM[0] = 128'h00C0006F063006132900081300000513;
      // RAM[1] = 128'h40B806B30025159302C50A6300150513;
      // RAM[2] = 128'hFED702E30047071300C0006F10400713;
      // RAM[3] = 128'hFEB72E23FEF5D8E300072583FFC72783;
      // RAM[4] = 128'h0000806700000513FE5FF06F00F72023;
  end


  always @(posedge clk)
    if (we)
      begin

        RAM[a[13:4]] <= wd;

  	  end
endmodule

/*
冒泡排序0-100，初始地址0x00000100
0x00000513
0x29000813
0x06300613
0x00C0006F

0x00150513
0x02C50A63
0x00251593
0x40B806B3

0x10400713
0x00C0006F
0x00470713
0xFED702E3

0xFFC72783
0x00072583
0xFEF5D8E3
0xFEB72E23

0x00F72023
0xFE5FF06F
0x00000513
0x00008067
*/